// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

////////////////////////////////////////////////////////////////////////////////
// Engineer:       Renzo Andri - andrire@student.ethz.ch                      //
//                                                                            //
// Additional contributions by:                                               //
//                 Igor Loi - igor.loi@unibo.it                               //
//                 Andreas Traber - atraber@student.ethz.ch                   //
//                 Sven Stucki - svstucki@student.ethz.ch                     //
//                                                                            //
// Design Name:    Instruction Fetch Stage                                    //
// Project Name:   RI5CY                                                      //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    Instruction fetch unit: Selection of the next PC, and      //
//                 buffering (sampling) of the read instruction               //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

module cv32e40p_if_stage #(
    parameter COREV_PULP = 0, // PULP ISA Extension (including PULP specific CSRs and hardware loop, excluding cv.elw)
    parameter PULP_OBI = 0,  // Legacy PULP OBI behavior
    parameter PULP_SECURE = 0,
    parameter FPU = 0,
    parameter ZFINX = 0
) (
    input logic clk,
    input logic rst_n,

    // Used to calculate the exception offsets
    input logic [23:0] m_trap_base_addr_i,
    input logic [23:0] u_trap_base_addr_i,
    input logic [ 1:0] trap_addr_mux_i,
    // Boot address
    input logic [31:0] boot_addr_i,
    input logic [31:0] dm_exception_addr_i,

    // Debug mode halt address
    input logic [31:0] dm_halt_addr_i,

    // instruction request control
    input logic req_i,

    // instruction cache interface
    output logic instr_req_o,
    output logic [31:0] instr_addr_o,
    input logic instr_gnt_i,
    input logic instr_rvalid_i,
    input logic [31:0] instr_rdata_i,
    input logic instr_err_i,      // External bus error (validity defined by instr_rvalid_i) (not used yet)
    input logic instr_err_pmp_i,  // PMP error (validity defined by instr_gnt_i)

    // Output of IF Pipeline stage
    output logic instr_valid_id_o,  // instruction in IF/ID pipeline is valid
    output logic [31:0] instr_rdata_id_o,      // read instruction is sampled and sent to ID stage for decoding
    output logic is_compressed_id_o,  // compressed decoder thinks this is a compressed instruction
    output logic illegal_c_insn_id_o,  // compressed decoder thinks this is an invalid instruction
    output logic [31:0] pc_if_o,
    output logic [31:0] pc_id_o,
    output logic is_fetch_failed_o,

    // Forwarding ports - control signals
    input logic clear_instr_valid_i,  // clear instruction valid bit in IF/ID pipe
    input logic pc_set_i,  // set the program counter to a new value
    input logic [31:0] mepc_i,  // address used to restore PC when the interrupt/exception is served
    input logic [31:0] uepc_i,  // address used to restore PC when the interrupt/exception is served

    input logic [31:0] depc_i,  // address used to restore PC when the debug is served

    input logic [3:0] pc_mux_i,  // sel for pc multiplexer
    input logic [2:0] exc_pc_mux_i,  // selects ISR address

    input  logic [4:0] m_exc_vec_pc_mux_i,  // selects ISR address for vectorized interrupt lines
    input  logic [4:0] u_exc_vec_pc_mux_i,  // selects ISR address for vectorized interrupt lines
    output logic       csr_mtvec_init_o,  // tell CS regfile to init mtvec

    // jump and branch target and decision
    input logic [31:0] jump_target_id_i,  // jump target address
    input logic [31:0] jump_target_ex_i,  // jump target address

    // from hwloop controller
    input logic        hwlp_jump_i,
    input logic [31:0] hwlp_target_i,

    // pipeline stall
    input logic halt_if_i,
    input logic id_ready_i,

    // misc signals
    output logic if_busy_o,  // is the IF stage busy fetching instructions?
    output logic perf_imiss_o,  // Instruction Fetch Miss
    //Error Detection Ports
    output logic error_detected_if1,
    output logic error_detected_if2,
    output logic error_detected_dec,
    output logic error_detected_dec2,
    output logic error_detected_dec3,
    output logic error_detected_dec4,
    output logic error_detected_dec5,
    output logic error_detected_dec6,
    output logic error_detected_dec7,
    output logic error_detected_dec8,
    
    output logic error_prefech_buffer_parity_o
);

  import cv32e40p_pkg::*;

  logic if_valid, if_ready;

  // prefetch buffer related signals
  logic        prefetch_busy;
  logic        branch_req;
  logic [31:0] branch_addr_n;
  logic [31:0] branch_addr_n2;

  logic        fetch_valid;
  logic        fetch_ready;
  logic [31:0] fetch_rdata;

  logic [31:0] exc_pc;
  logic [31:0] exc_pc2;

  logic [23:0] trap_base_addr;
  logic [ 4:0] exc_vec_pc_mux;
  logic        fetch_failed;

  logic        aligner_ready;
  logic        instr_valid;

  logic        illegal_c_insn;
  logic [31:0] instr_aligned;
  logic [31:0] instr_decompressed;
  logic        instr_compressed_int;


  // exception PC selection mux
  always_comb begin : EXC_PC_MUX
    unique case (trap_addr_mux_i)
      TRAP_MACHINE: trap_base_addr = m_trap_base_addr_i;
      TRAP_USER:    trap_base_addr = u_trap_base_addr_i;
      default:      trap_base_addr = m_trap_base_addr_i;
    endcase

    unique case (trap_addr_mux_i)
      TRAP_MACHINE: exc_vec_pc_mux = m_exc_vec_pc_mux_i;
      TRAP_USER:    exc_vec_pc_mux = u_exc_vec_pc_mux_i;
      default:      exc_vec_pc_mux = m_exc_vec_pc_mux_i;
    endcase

    unique case (exc_pc_mux_i)
      EXC_PC_EXCEPTION:
      exc_pc = {trap_base_addr, 8'h0};  //1.10 all the exceptions go to base address
      EXC_PC_IRQ: exc_pc = {trap_base_addr, 1'b0, exc_vec_pc_mux, 2'b0};  // interrupts are vectored
      EXC_PC_DBD: exc_pc = {dm_halt_addr_i[31:2], 2'b0};
      EXC_PC_DBE: exc_pc = {dm_exception_addr_i[31:2], 2'b0};
      default: exc_pc = {trap_base_addr, 8'h0};
    endcase
    unique case (exc_pc_mux_i)
      EXC_PC_EXCEPTION:
      exc_pc2 = {trap_base_addr, 8'h0};  //1.10 all the exceptions go to base address
      EXC_PC_IRQ: exc_pc2 = {trap_base_addr, 1'b0, exc_vec_pc_mux, 2'b0};  // interrupts are vectored
      EXC_PC_DBD: exc_pc2 = {dm_halt_addr_i[31:2], 2'b0};
      EXC_PC_DBE: exc_pc2 = {dm_exception_addr_i[31:2], 2'b0};
      default: exc_pc2 = {trap_base_addr, 8'h0};
    endcase

    if (exc_pc != exc_pc2) begin
      error_detected_if1 = 1;
    end else begin
      error_detected_if1 = 0;
    end
  end

  // fetch address selection
  always_comb begin
    // Default assign PC_BOOT (should be overwritten in below case)
    branch_addr_n = {boot_addr_i[31:2], 2'b0};
    branch_addr_n2 = {boot_addr_i[31:2], 2'b0};

    unique case (pc_mux_i)
      PC_BOOT: branch_addr_n = {boot_addr_i[31:2], 2'b0};
      PC_JUMP: branch_addr_n = jump_target_id_i;
      PC_BRANCH: branch_addr_n = jump_target_ex_i;
      PC_EXCEPTION: branch_addr_n = exc_pc;  // set PC to exception handler
      PC_MRET: branch_addr_n = mepc_i;  // PC is restored when returning from IRQ/exception
      PC_URET: branch_addr_n = uepc_i;  // PC is restored when returning from IRQ/exception
      PC_DRET: branch_addr_n = depc_i;  //
      PC_FENCEI: branch_addr_n = pc_id_o + 4;  // jump to next instr forces prefetch buffer reload
      PC_HWLOOP: branch_addr_n = hwlp_target_i;
      default: ;
    endcase
    unique case (pc_mux_i)
      PC_BOOT: branch_addr_n2 = {boot_addr_i[31:2], 2'b0};
      PC_JUMP: branch_addr_n2 = jump_target_id_i;
      PC_BRANCH: branch_addr_n2 = jump_target_ex_i;
      PC_EXCEPTION: branch_addr_n2 = exc_pc;  // set PC to exception handler
      PC_MRET: branch_addr_n2 = mepc_i;  // PC is restored when returning from IRQ/exception
      PC_URET: branch_addr_n2 = uepc_i;  // PC is restored when returning from IRQ/exception
      PC_DRET: branch_addr_n2 = depc_i;  //
      PC_FENCEI: branch_addr_n2 = pc_id_o + 4;  // jump to next instr forces prefetch buffer reload
      PC_HWLOOP: branch_addr_n2 = hwlp_target_i;
      default: ;
    endcase

    if(branch_addr_n != branch_addr_n2) begin
      error_detected_if2 = 1;
    end else begin
      error_detected_if2 = 0;
    end
  end

  // tell CS register file to initialize mtvec on boot
  assign csr_mtvec_init_o = (pc_mux_i == PC_BOOT) & pc_set_i;

  assign fetch_failed    = 1'b0; // PMP is not supported in CV32E40P

  // prefetch buffer, caches a fixed number of instructions
  cv32e40p_prefetch_buffer #(
      .PULP_OBI  (PULP_OBI),
      .COREV_PULP(COREV_PULP)
  ) prefetch_buffer_i (
      .clk  (clk),
      .rst_n(rst_n),

      .req_i(req_i),

      .branch_i     (branch_req),
      .branch_addr_i({branch_addr_n[31:1], 1'b0}),

      .hwlp_jump_i  (hwlp_jump_i),
      .hwlp_target_i(hwlp_target_i),

      .fetch_ready_i(fetch_ready),
      .fetch_valid_o(fetch_valid),
      .fetch_rdata_o(fetch_rdata),

      // goes to instruction memory / instruction cache
      .instr_req_o    (instr_req_o),
      .instr_addr_o   (instr_addr_o),
      .instr_gnt_i    (instr_gnt_i),
      .instr_rvalid_i (instr_rvalid_i),
      .instr_err_i    (instr_err_i),  // Not supported (yet)
      .instr_err_pmp_i(instr_err_pmp_i),  // Not supported (yet)
      .instr_rdata_i  (instr_rdata_i),

      // Prefetch Buffer Status
      .busy_o(prefetch_busy),

      .error_prefech_buffer_parity_o(error_prefech_buffer_parity_o)
  );

  // offset FSM state transition logic
  always_comb begin

    fetch_ready = 1'b0;
    branch_req  = 1'b0;
    // take care of jumps and branches
    if (pc_set_i) begin
      branch_req = 1'b1;
    end else if (fetch_valid) begin
      if (req_i && if_valid) begin
        fetch_ready = aligner_ready;
      end
    end
  end

  assign if_busy_o    = prefetch_busy;
  assign perf_imiss_o = !fetch_valid && !branch_req;

  // IF-ID pipeline registers, frozen when the ID stage is stalled
  always_ff @(posedge clk, negedge rst_n) begin : IF_ID_PIPE_REGISTERS
    if (rst_n == 1'b0) begin
      instr_valid_id_o    <= 1'b0;
      instr_rdata_id_o    <= '0;
      is_fetch_failed_o   <= 1'b0;
      pc_id_o             <= '0;
      is_compressed_id_o  <= 1'b0;
      illegal_c_insn_id_o <= 1'b0;
    end else begin

      if (if_valid && instr_valid) begin
        instr_valid_id_o    <= 1'b1;
        instr_rdata_id_o    <= instr_decompressed;
        is_compressed_id_o  <= instr_compressed_int;
        illegal_c_insn_id_o <= illegal_c_insn;
        is_fetch_failed_o   <= 1'b0;
        pc_id_o             <= pc_if_o;
      end else if (clear_instr_valid_i) begin
        instr_valid_id_o  <= 1'b0;
        is_fetch_failed_o <= fetch_failed;
      end
    end
  end

  assign if_ready = fetch_valid & id_ready_i;
  assign if_valid = (~halt_if_i) & if_ready;

  cv32e40p_aligner aligner_i (
      .clk             (clk),
      .rst_n           (rst_n),
      .fetch_valid_i   (fetch_valid),
      .aligner_ready_o (aligner_ready),
      .if_valid_i      (if_valid),
      .fetch_rdata_i   (fetch_rdata),
      .instr_aligned_o (instr_aligned),
      .instr_valid_o   (instr_valid),
      .branch_addr_i   ({branch_addr_n[31:1], 1'b0}),
      .branch_i        (branch_req),
      .hwlp_addr_i     (hwlp_target_i),
      .hwlp_update_pc_i(hwlp_jump_i),
      .pc_o            (pc_if_o)
  );


  logic [31:0] instr_decompressed1;
  logic [31:0] instr_decompressed_mux1, instr_decompressed_mux2;

  cv32e40p_compressed_decoder #(
      .FPU  (FPU),
      .ZFINX(ZFINX)
  ) compressed_decoder_i (
      .instr_i        (instr_aligned),
      .instr_o        (instr_decompressed1),
      .is_compressed_o(instr_compressed_int),
      .illegal_instr_o(illegal_c_insn)
  );

  logic [31:0] instr_decompressed2;

  cv32e40p_compressed_decoder #(
      .FPU  (FPU),
      .ZFINX(ZFINX)
  ) compressed_decoder_i2 (
      .instr_i        (instr_aligned),
      .instr_o        (instr_decompressed2),
      .is_compressed_o(instr_compressed_int2),
      .illegal_instr_o(illegal_c_insn2)
  );


  logic [31:0] instr_decompressed3;

  cv32e40p_compressed_decoder #(
      .FPU  (FPU),
      .ZFINX(ZFINX)
  ) compressed_decoder_i3 (
      .instr_i        (instr_aligned),
      .instr_o        (instr_decompressed3),
      .is_compressed_o(instr_compressed_int3),
      .illegal_instr_o(illegal_c_insn3)
  );

  logic [31:0] instr_decompressed4;

  cv32e40p_compressed_decoder #(
      .FPU  (FPU),
      .ZFINX(ZFINX)
  ) compressed_decoder_i4 (
      .instr_i        (instr_aligned),
      .instr_o        (instr_decompressed4),
      .is_compressed_o(instr_compressed_int4),
      .illegal_instr_o(illegal_c_insn4)
  );

  logic [31:0] instr_decompressed5;

  cv32e40p_compressed_decoder #(
      .FPU  (FPU),
      .ZFINX(ZFINX)
  ) compressed_decoder_i5 (
      .instr_i        (instr_aligned),
      .instr_o        (instr_decompressed5),
      .is_compressed_o(instr_compressed_int5),
      .illegal_instr_o(illegal_c_insn5)
  );

  logic [31:0] instr_decompressed6;

  cv32e40p_compressed_decoder #(
      .FPU  (FPU),
      .ZFINX(ZFINX)
  ) compressed_decoder_i6 (
      .instr_i        (instr_aligned),
      .instr_o        (instr_decompressed6),
      .is_compressed_o(instr_compressed_int),
      .illegal_instr_o(illegal_c_insn)
  );

  logic [31:0] instr_decompressed7;

  cv32e40p_compressed_decoder #(
      .FPU  (FPU),
      .ZFINX(ZFINX)
  ) compressed_decoder_i7 (
      .instr_i        (instr_aligned),
      .instr_o        (instr_decompressed7),
      .is_compressed_o(instr_compressed_int),
      .illegal_instr_o(illegal_c_insn)
  );

  logic [31:0] instr_decompressed8;

  cv32e40p_compressed_decoder #(
      .FPU  (FPU),
      .ZFINX(ZFINX)
  ) compressed_decoder_i8 (
      .instr_i        (instr_aligned),
      .instr_o        (instr_decompressed8),
      .is_compressed_o(instr_compressed_int),
      .illegal_instr_o(illegal_c_insn)
  );

  logic [31:0] instr_decompressed9;

  cv32e40p_compressed_decoder #(
      .FPU  (FPU),
      .ZFINX(ZFINX)
  ) compressed_decoder_i9 (
      .instr_i        (instr_aligned),
      .instr_o        (instr_decompressed9),
      .is_compressed_o(instr_compressed_int),
      .illegal_instr_o(illegal_c_insn)
  );

  logic [1:0] selMUX;
  logic selMUX_o;

  always_comb begin
    
    if (instr_decompressed1 != instr_decompressed2) begin
      error_detected_dec = 1;
    end else begin
      error_detected_dec = 0;
    end
    if (instr_decompressed1 != instr_decompressed3) begin
        error_detected_dec2 = 1;
    end else begin
      error_detected_dec2 = 0;
    end
  
    if (instr_decompressed1 != instr_decompressed4) begin
        error_detected_dec3 = 1;
    end else begin
      error_detected_dec3 = 0;
    end

    if (instr_decompressed1 != instr_decompressed5) begin
        error_detected_dec4 = 1;
    end else begin
      error_detected_dec4 = 0;
    end

    if (instr_decompressed1 != instr_decompressed6) begin
      error_detected_dec5 = 1;
    end else begin
      error_detected_dec5 = 0;
    end
    if (instr_decompressed1 != instr_decompressed7) begin
        error_detected_dec6 = 1;
    end else begin
      error_detected_dec6 = 0;
    end
  
    if (instr_decompressed1 != instr_decompressed8) begin
        error_detected_dec7 = 1;
    end else begin
      error_detected_dec7 = 0;
    end

    if (instr_decompressed9 != instr_decompressed9) begin
        error_detected_dec8 = 1;
    end else begin
      error_detected_dec8 = 0;
    end


    selMUX[1] = error_detected_dec & error_detected_dec2;
    selMUX[0] = (error_detected_dec & ~error_detected_dec2) | (error_detected_dec & error_detected_dec2 & error_detected_dec3);
    selMUX_o = error_detected_dec & error_detected_dec2 & error_detected_dec3 & error_detected_dec4 ;
    //selMUX_mult = error_detected_mult & ~error_detected_mult2;

    //the MUX implementation
    
    case(selMUX)

	      2'b00: begin instr_decompressed_mux1 = instr_decompressed1; end
        2'b01: begin instr_decompressed_mux1 = instr_decompressed2; end
        2'b10: begin instr_decompressed_mux1 = instr_decompressed3; end
        default: begin instr_decompressed_mux1 = instr_decompressed4; end

    endcase

    case(selMUX)

	      2'b00: begin instr_decompressed_mux2 = instr_decompressed5; end
        2'b01: begin instr_decompressed_mux2 = instr_decompressed6; end
        2'b10: begin instr_decompressed_mux2 = instr_decompressed7; end
        default: begin instr_decompressed_mux2 = instr_decompressed8; end

    endcase

    case(selMUX_o)

        1'b0: begin instr_decompressed = instr_decompressed_mux1; end
        default: begin instr_decompressed = instr_decompressed_mux2; end

    endcase

  end
  //----------------------------------------------------------------------------
  // Assertions
  //----------------------------------------------------------------------------

`ifdef CV32E40P_ASSERT_ON

  generate
    if (!COREV_PULP) begin : gen_no_pulp_xpulp_assertions

      // Check that PC Mux cannot select Hardware Loop address iF PULP extensions are not included
      property p_pc_mux_0;
        @(posedge clk) disable iff (!rst_n) (1'b1) |-> (pc_mux_i != PC_HWLOOP);
      endproperty

      a_pc_mux_0 :
      assert property (p_pc_mux_0);

    end
  endgenerate

  generate
    if (!PULP_SECURE) begin : gen_no_pulp_secure_assertions

      // Check that PC Mux cannot select URET address if User Mode is not included
      property p_pc_mux_1;
        @(posedge clk) disable iff (!rst_n) (1'b1) |-> (pc_mux_i != PC_URET);
      endproperty

      a_pc_mux_1 :
      assert property (p_pc_mux_1);

    end
  endgenerate

`endif

endmodule

// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// Top file instantiating a CV32E40P core and an optional FPU
// Contributor: Davide Schiavone <davide@openhwgroup.org>

module cv32e40p_top #(
    parameter COREV_PULP = 0, // PULP ISA Extension (incl. custom CSRs and hardware loop, excl. cv.elw)
    parameter COREV_CLUSTER = 0,  // PULP Cluster interface (incl. cv.elw)
    parameter FPU = 0,  // Floating Point Unit (interfaced via APU interface)
    parameter FPU_ADDMUL_LAT = 0,  // Floating-Point ADDition/MULtiplication computing lane pipeline registers number
    parameter FPU_OTHERS_LAT = 0,  // Floating-Point COMParison/CONVersion computing lanes pipeline registers number
    parameter ZFINX = 0,  // Float-in-General Purpose registers
    parameter NUM_MHPMCOUNTERS = 1
) (
    // Clock and Reset
    input logic clk_i,
    input logic rst_ni,

    input logic pulp_clock_en_i,  // PULP clock enable (only used if COREV_CLUSTER = 1)
    input logic scan_cg_en_i,  // Enable all clock gates for testing

    // Core ID, Cluster ID, debug mode halt address and boot address are considered more or less static
    input logic [31:0] boot_addr_i,
    input logic [31:0] mtvec_addr_i,
    input logic [31:0] dm_halt_addr_i,
    input logic [31:0] hart_id_i,
    input logic [31:0] dm_exception_addr_i,

    // Instruction memory interface
    output logic        instr_req_o,
    input  logic        instr_gnt_i,
    input  logic        instr_rvalid_i,
    output logic [31:0] instr_addr_o,
    input  logic [31:0] instr_rdata_i,

    // Data memory interface
    output logic        data_req_o,
    input  logic        data_gnt_i,
    input  logic        data_rvalid_i,
    output logic        data_we_o,
    output logic [ 3:0] data_be_o,
    output logic [31:0] data_addr_o,
    output logic [31:0] data_wdata_o,
    input  logic [31:0] data_rdata_i,

    // Interrupt inputs
    input  logic [31:0] irq_i,  // CLINT interrupts + CLINT extension interrupts
    output logic        irq_ack_o,
    output logic [ 4:0] irq_id_o,

    // Debug Interface
    input  logic debug_req_i,
    output logic debug_havereset_o,
    output logic debug_running_o,
    output logic debug_halted_o,

    // CPU Control Signals
    input  logic fetch_enable_i,
    output logic core_sleep_o,
    //Error Detection Ports
    output logic error_detected_ex1,
    output logic error_detected_alu,
    output logic error_detected_alu2,
    output logic error_detected_alu3,
    output logic error_detected_alu4,
    output logic error_detected_alu5,
    output logic error_detected_alu6,
    output logic error_detected_alu7,
    output logic error_detected_alu8,
    output logic error_detected_mult,
    output logic error_detected_mult2,
    output logic error_detected_mult3,
    output logic error_detected_mult4,
    output logic error_detected_mult5,
    output logic error_detected_mult6,
    output logic error_detected_mult7,
    output logic error_detected_mult8,
    output logic error_detected_if1,
    output logic error_detected_if2,
    output logic error_detected_dec,
    output logic error_detected_dec2,
    output logic error_detected_dec3,
    output logic error_detected_dec4,
    output logic error_detected_dec5,
    output logic error_detected_dec6,
    output logic error_detected_dec7,
    output logic error_detected_dec8,
    output logic error_detected_id1,
    output logic error_detected_id2,
    output logic error_detected_id3,

    output logic [5:0]			error_parity_regfile_o,
	  //output logic [3:0]			error_decoder_o,
	  output logic [2:0]			error_parity_id_ex_stage_o,
	  output logic [3:0]			error_load_store_o,
	  output logic 				error_prefech_buffer_parity_o,

    output logic error_detected_decod1,
    output logic error_detected_decod2,
    output logic error_detected_decod3
);

  import cv32e40p_apu_core_pkg::*;

  // Core to FPU
  logic                              clk;
  logic                              apu_req;
  logic [   APU_NARGS_CPU-1:0][31:0] apu_operands;
  logic [     APU_WOP_CPU-1:0]       apu_op;
  logic [APU_NDSFLAGS_CPU-1:0]       apu_flags;

  // FPU to Core
  logic                              apu_gnt;
  logic                              apu_rvalid;
  logic [                31:0]       apu_rdata;
  logic [APU_NUSFLAGS_CPU-1:0]       apu_rflags;

  // Instantiate the Core
  cv32e40p_core #(
      .COREV_PULP      (COREV_PULP),
      .COREV_CLUSTER   (COREV_CLUSTER),
      .FPU             (FPU),
      .FPU_ADDMUL_LAT  (FPU_ADDMUL_LAT),
      .FPU_OTHERS_LAT  (FPU_OTHERS_LAT),
      .ZFINX           (ZFINX),
      .NUM_MHPMCOUNTERS(NUM_MHPMCOUNTERS)
  ) core_i (
      .clk_i (clk_i),
      .rst_ni(rst_ni),

      .pulp_clock_en_i(pulp_clock_en_i),
      .scan_cg_en_i   (scan_cg_en_i),

      .boot_addr_i        (boot_addr_i),
      .mtvec_addr_i       (mtvec_addr_i),
      .dm_halt_addr_i     (dm_halt_addr_i),
      .hart_id_i          (hart_id_i),
      .dm_exception_addr_i(dm_exception_addr_i),

      .instr_req_o   (instr_req_o),
      .instr_gnt_i   (instr_gnt_i),
      .instr_rvalid_i(instr_rvalid_i),
      .instr_addr_o  (instr_addr_o),
      .instr_rdata_i (instr_rdata_i),

      .data_req_o   (data_req_o),
      .data_gnt_i   (data_gnt_i),
      .data_rvalid_i(data_rvalid_i),
      .data_we_o    (data_we_o),
      .data_be_o    (data_be_o),
      .data_addr_o  (data_addr_o),
      .data_wdata_o (data_wdata_o),
      .data_rdata_i (data_rdata_i),

      .apu_req_o     (apu_req),
      .apu_gnt_i     (apu_gnt),
      .apu_operands_o(apu_operands),
      .apu_op_o      (apu_op),
      .apu_flags_o   (apu_flags),
      .apu_rvalid_i  (apu_rvalid),
      .apu_result_i  (apu_rdata),
      .apu_flags_i   (apu_rflags),

      .irq_i    (irq_i),
      .irq_ack_o(irq_ack_o),
      .irq_id_o (irq_id_o),

      .debug_req_i      (debug_req_i),
      .debug_havereset_o(debug_havereset_o),
      .debug_running_o  (debug_running_o),
      .debug_halted_o   (debug_halted_o),

      .fetch_enable_i(fetch_enable_i),
      .core_sleep_o  (core_sleep_o),
      
      .error_detected_ex1(error_detected_ex1),
      .error_detected_alu (error_detected_alu),
      .error_detected_alu2 (error_detected_alu2),
      .error_detected_alu3(error_detected_alu3),
      .error_detected_alu4(error_detected_alu4),
      .error_detected_alu5(error_detected_alu5),
      .error_detected_alu6(error_detected_alu6),
      .error_detected_alu7(error_detected_alu7),
      .error_detected_alu8(error_detected_alu8),
      .error_detected_mult(error_detected_mult),
      .error_detected_mult2(error_detected_mult2),
      .error_detected_mult3(error_detected_mult3),
      .error_detected_mult4(error_detected_mult4),
      .error_detected_mult5(error_detected_mult5),
      .error_detected_mult6(error_detected_mult6),
      .error_detected_mult7(error_detected_mult7),
      .error_detected_mult8(error_detected_mult8),
      .error_detected_if1(error_detected_if1),
      .error_detected_if2(error_detected_if2),
      .error_detected_dec(error_detected_dec),
      .error_detected_dec2(error_detected_dec2),
      .error_detected_dec3(error_detected_dec3),
      .error_detected_dec4(error_detected_dec4),
      .error_detected_dec5(error_detected_dec5),
      .error_detected_dec6(error_detected_dec6),
      .error_detected_dec7(error_detected_dec7),
      .error_detected_dec8(error_detected_dec8),
      .error_detected_id1(error_detected_id1),
      .error_detected_id2(error_detected_id2),
      .error_detected_id3(error_detected_id3),

      .error_parity_regfile_o(error_parity_regfile_o),
	    //.error_decoder_o(error_decoder_o),
	    .error_parity_id_ex_stage_o(error_parity_id_ex_stage_o),
	    .error_load_store_o(error_load_store_o),
	    .error_prefech_buffer_parity_o(error_prefech_buffer_parity_o),

      .error_detected_decod1(error_detected_decod1),
      .error_detected_decod2(error_detected_decod2),
      .error_detected_decod3(error_detected_decod3)
  );

  generate
    if (FPU) begin : fpu_gen
      // FPU clock gate
      cv32e40p_clock_gate core_clock_gate_i (
          .clk_i       (clk_i),
          .en_i        (!core_sleep_o),
          .scan_cg_en_i(scan_cg_en_i),
          .clk_o       (clk)
      );

      // Instantiate the FPU wrapper
      cv32e40p_fp_wrapper #(
          .FPU_ADDMUL_LAT(FPU_ADDMUL_LAT),
          .FPU_OTHERS_LAT(FPU_OTHERS_LAT)
      ) fp_wrapper_i (
          .clk_i         (clk),
          .rst_ni        (rst_ni),
          .apu_req_i     (apu_req),
          .apu_gnt_o     (apu_gnt),
          .apu_operands_i(apu_operands),
          .apu_op_i      (apu_op),
          .apu_flags_i   (apu_flags),
          .apu_rvalid_o  (apu_rvalid),
          .apu_rdata_o   (apu_rdata),
          .apu_rflags_o  (apu_rflags)
      );
    end else begin : no_fpu_gen
      // Drive FPU output signals to 0
      assign apu_gnt    = '0;
      assign apu_rvalid = '0;
      assign apu_rdata  = '0;
      assign apu_rflags = '0;
    end
  endgenerate

endmodule
